module example_top (
    input a,
    input b,

    output c
);

or_gate or_gate_top (
    .a,
    .b,
    .c
);

endmodule
